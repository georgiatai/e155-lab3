/////////////////////////
// lab3_gt.sv
// Author: Georgia Tai, ytai@g.hmc.edu
// Date: Sep 14, 2025
// 
// Top level module for Lab 3 of E155 @HMC. 
// Takes in a 4-by-4 keypad and uses dual seven segment display to 
// show the most recent two inputs.
/////////////////////////

